`include "defines.v"
module mips(
	input wire	clk,
	input wire	rst,

	input wire[`RegBus]	rom_data_i,
	input wire[`RegBus]	ram_data_i,
	
	output wire[`RegBus]	rom_addr_o,
	output wire		rom_ce_o,

	output wire[`RegBus]	ram_addr_o,
	output wire[`RegBus]	ram_data_o,
	output wire		ram_we_o,
	output wire[3:0]	ram_sel_o,
	output wire		ram_ce_o
);

// connect IF/ID with ID
wire[`InstAddrBus] 	pc;
wire[`InstAddrBus] 	id_pc_i;
wire[`InstBus] 		id_inst_i;

//connect ID with ID/EX
wire[`AluOpBus]		id_aluop_o;
wire[`AluSelBus]	id_alusel_o;
wire[`RegBus]		id_reg1_o;
wire[`RegBus]		id_reg2_o;
wire			id_wreg_o;
wire[`RegAddrBus]	id_wd_o;

//connect ID/EX with EX
wire[`AluOpBus]		ex_aluop_i;
wire[`AluSelBus] 	ex_alusel_i;
wire[`RegBus] 		ex_reg1_i;
wire[`RegBus]		ex_reg2_i;
wire			ex_wreg_i;
wire[`RegAddrBus]	ex_wd_i;

//connect EX with EX/MEM
wire 			ex_wreg_o;
wire[`RegAddrBus]	ex_wd_o;
wire[`RegBus]		ex_wdata_o;

//connect EX/MEM with MEM
wire 			mem_wreg_i;
wire[`RegAddrBus]	mem_wd_i;
wire[`RegBus]		mem_wdata_i;

//connect MEM with MEM/WB
wire 			mem_wreg_o;
wire[`RegAddrBus]	mem_wd_o;
wire[`RegBus]		mem_wdata_o;

//connect MEM/wb with wb
wire 			wb_wreg_i;
wire[`RegAddrBus]	wb_wd_i;
wire[`RegBus]		wb_wdata_i;

// connect ID with RegFile
wire 			reg1_read;
wire			reg2_read;
wire[`RegBus]		reg1_data;
wire[`RegBus]		reg2_data;
wire[`RegAddrBus]	reg1_addr;
wire[`RegAddrBus]	reg2_addr;

// about branch
// IN ID
wire[`RegBus] 		id_branch_target_address_o;
wire 			id_branch_flag_o;
wire			id_next_inst_in_delayslot_o;
wire[`RegBus]		id_link_addr_o;
wire			id_is_in_delayslot_o;

// IN ID/EX
wire[`RegBus]		ex_link_address;
wire			ex_is_in_delayslot;
wire			ex_is_in_delayslot_o;

//memory
wire[`InstBus]		id_ex_inst;
wire[`InstBus]		ex_inst;

wire[`AluOpBus]		ex_aluop_o;
wire[`RegBus]		ex_mem_addr_o;
wire[`RegBus]		ex_reg2_o;
wire[`AluOpBus]		mem_aluop_o;
wire[`RegBus]		mem_mem_addr_o;
wire[`RegBus]		mem_reg2_o;

//control
wire[5:0]		stall;
wire			stallreq_from_id;
wire			stallreq_from_ex;

//instance PC
pc U_PC (
	.clk(clk), .rst(rst),.pc(pc),
	.ce(rom_ce_o),.stall(stall),
	.branch_flag_i(id_branch_flag_o),.branch_target_address_i(id_branch_target_address_o)
);

assign rom_addr_o = pc;		//the address of ROM INPUT == PC

// instance IF/ID
if_id U_IF_ID (
	.clk(clk), .rst(rst), .if_pc(pc),.stall(stall),
	.if_inst(rom_data_i),.id_pc(id_pc_i),
	.id_inst(id_inst_i)
);

//instance ID
id U_ID (
	.rst(rst), .pc_i(id_pc_i),.inst_i(id_inst_i),
	// from RegFile
	.reg1_data_i(reg1_data), .reg2_data_i(reg2_data),
	
	//from EX to avoid RAW
	.ex_wreg_i(ex_wreg_o),.ex_wdata_i(ex_wdata_o),
	.ex_wd_i(ex_wd_o),

	//from EX to avoid Load About
	.ex_aluop_i(ex_aluop_o),	

	//from MEM to avoid RAW
	.mem_wreg_i(mem_wreg_o),.mem_wdata_i(mem_wdata_o),
	.mem_wd_i(mem_wd_o),

	// to RegFile
	.reg1_read_o(reg1_read),.reg2_read_o(reg2_read),
	.reg1_addr_o(reg1_addr),.reg2_addr_o(reg2_addr),
	
	//branch
	.is_in_delayslot_i(ex_is_in_delayslot_o),

	.branch_flag_o(id_branch_flag_o),.branch_target_address_o(id_branch_target_address_o),
	.next_inst_in_delayslot_o(id_next_inst_in_delayslot_o),.is_in_delayslot_o(id_is_in_delayslot_o),
	.link_addr_o(id_link_addr_o),

	// to ID/EX
	.aluop_o(id_aluop_o),.alusel_o(id_alusel_o),
	.reg1_o(id_reg1_o),.reg2_o(id_reg2_o),
	.wd_o(id_wd_o),.wreg_o(id_wreg_o),

	//memory
	.inst_o(id_ex_inst),
	
	//to control
	.stallreq(stallreq_from_id)
);

//instance RegFile
regfile U_REGFILE(
	.clk(clk),	.rst(rst),
	.we(wb_wreg_i),	.waddr(wb_wd_i),
	.wdata(wb_wdata_i),
	.re1(reg1_read),
	.raddr1(reg1_addr),.rdata1(reg1_data),
	.re2(reg2_read),
	.raddr2(reg2_addr),.rdata2(reg2_data)
);

//instance ID/EX
id_ex U_ID_EX (
	.clk(clk),	.rst(rst),	.stall(stall),
	
	.id_aluop(id_aluop_o),	.id_alusel(id_alusel_o),
	.id_reg1(id_reg1_o),	.id_reg2(id_reg2_o),
	.id_wd(id_wd_o),	.id_wreg(id_wreg_o),
	.id_is_in_delayslot(id_is_in_delayslot_o),	.id_link_address(id_link_addr_o),
	.next_inst_in_delayslot_i(id_next_inst_in_delayslot_o),	

	.ex_aluop(ex_aluop_i),	.ex_alusel(ex_alusel_i),
	.ex_reg1(ex_reg1_i),	.ex_reg2(ex_reg2_i),
	.ex_wd(ex_wd_i),	.ex_wreg(ex_wreg_i),
	.ex_is_in_delayslot(ex_is_in_delayslot),	.ex_link_address(ex_link_address),
	.is_in_delayslot_o(ex_is_in_delayslot_o),

	.id_inst(id_ex_inst),.ex_inst(ex_inst)

);

//instance ex
ex U_EX(
	.rst(rst),
	
	.aluop_i(ex_aluop_i),	.alusel_i(ex_alusel_i),
	.reg1_i(ex_reg1_i),	.reg2_i(ex_reg2_i),
	.wd_i(ex_wd_i),		.wreg_i(ex_wreg_i),
	.is_in_delayslot_i(ex_is_in_delayslot),	.link_address_i(ex_link_address),

	.wd_o(ex_wd_o),		.wreg_o(ex_wreg_o),
	.wdata_o(ex_wdata_o),
	
	.inst_i(ex_inst),.aluop_o(ex_aluop_o),
	.mem_addr_o(ex_mem_addr_o),.reg2_o(ex_reg2_o),

	//to control
	.stallreq(stallreq_from_ex)
);

ex_mem U_EX_MEM(
	.clk(clk),	.rst(rst),	.stall(stall),
	
	.ex_wd(ex_wd_o),		.ex_wreg(ex_wreg_o),
	.ex_wdata(ex_wdata_o),

	.mem_wd(mem_wd_i),		.mem_wreg(mem_wreg_i),
	.mem_wdata(mem_wdata_i),
	
	.ex_aluop(ex_aluop_o),		.ex_mem_addr(ex_mem_addr_o),
	.ex_reg2(ex_reg2_o),

	.mem_aluop(mem_aluop_o),.mem_mem_addr(mem_mem_addr_o),
	.mem_reg2(mem_reg2_o)
);

mem U_MEM(
	.rst(rst),
	.wd_i(mem_wd_i),		.wreg_i(mem_wreg_i),
	.wdata_i(mem_wdata_i),
	
	.aluop_i(mem_aluop_o),.mem_addr_i(mem_mem_addr_o),
	.reg2_i(mem_reg2_o),

	.mem_data_i(ram_data_i),	

	.wd_o(mem_wd_o),		.wreg_o(mem_wreg_o),
	.wdata_o(mem_wdata_o),

	.mem_addr_o(ram_addr_o),	.mem_we_o(ram_we_o),
	.mem_sel_o(ram_sel_o),		.mem_data_o(ram_data_o),
	.mem_ce_o(ram_ce_o)
);

mem_wb U_MEM_WB(
	.clk(clk),	.rst(rst),	.stall(stall),

	.mem_wd(mem_wd_o),		.mem_wreg(mem_wreg_o),
	.mem_wdata(mem_wdata_o),

	.wb_wd(wb_wd_i),		.wb_wreg(wb_wreg_i),
	.wb_wdata(wb_wdata_i)
);

control U_CONTROL(
	.rst(rst),
	.stallreq_from_id(stallreq_from_id),
	.stallreq_from_ex(stallreq_from_ex),
	.stall(stall)
);
endmodule