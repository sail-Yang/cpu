
`include "defines.v"
module mips_sopc(
	input wire	clk,
	input wire	rst
);

wire[`InstAddrBus]	inst_addr;
wire[`InstBus]		inst;

wire[`DataAddrBus]	data_addr;
wire[`DataBus]		data;
wire[`DataBus]		ram_data_o;
wire			rom_ce;
wire			ram_we;
wire			ram_ce;
wire[3:0]		ram_sel;

mips U_MIPS(
	.clk(clk),	.rst(rst),
	.rom_data_i(inst),.ram_data_i(data),
	.rom_addr_o(inst_addr), 
	.rom_ce_o(rom_ce),
	
	.ram_addr_o(data_addr),
	.ram_data_o(ram_data_o),
	.ram_we_o(ram_we),
	.ram_sel_o(ram_sel),
	.ram_ce_o(ram_ce)
);

im U_IM (
	.ce(rom_ce),
	.addr(inst_addr),
	.inst(inst)
);

dm U_DM (
	.clk(clk),.ce(ram_ce),.we(ram_we),
	.addr(data_addr),
	.sel(ram_sel),
	.data_i(ram_data_o),

	.data_o(data)
);

endmodule