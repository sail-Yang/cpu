
`include "defines.v"
module pc(
	input  wire			clk,
	input  wire			rst,
	
	input wire[5:0]			stall,
	//from module ID
	input wire			branch_flag_i,
	input wire[`RegBus]		branch_target_address_i,

	output reg[`InstAddrBus]	pc,
	output reg			ce

	
);

	always @ (posedge clk) begin
		if (rst == `RstEnable) begin
			ce <= `ChipDisable;	//When Reset,PC Disable
		end
		else begin
			ce <= `ChipEnable;
		end
	end
	
	always @ (posedge clk) begin
		if (ce == `ChipDisable) begin
			pc <= `InitAddr;	//When Disable,PC = 32'h00003000
		end else if(stall[0] == `NoStop) begin
			if(branch_flag_i == `Branch) begin
				pc <= branch_target_address_i;
			end else begin
				pc <= pc + 4'h4;	//pc += 4B,per clk 
			end
		end
	end
endmodule